// lab2.sv
// Description:
// Braden Vanderwoerd, 1/18/2026

module lab2_tb;

endmodule